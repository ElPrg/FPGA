   input    hsma_clk_in0_d_40_D_CLK,
   
   
	inout 	hsma_io_41_DATA0     , hsma_io_42_DATA16   ,
			hsma_io_43_DATA1     , hsma_io_44_DATA17   ,
			hsma_io_47_DATA2     , hsma_io_48_DATA18   ,
			hsma_io_49_DATA3     , hsma_io_50_DATA19   ,
			hsma_io_53_DATA4     , hsma_io_54_DATA20   ,
			hsma_io_55_DATA5     , hsma_io_56_DATA21   ,
			hsma_io_59_DATA6     , hsma_io_60_DATA22   ,
			hsma_io_61_DATA7     , hsma_io_62_DATA23   ,
			hsma_io_65_DATA8     , hsma_io_66_DATA24   ,
			hsma_io_67_DATA9     , hsma_io_68_DATA25   ,
			hsma_io_71_DATA10    , hsma_io_72_DATA26   ,
			hsma_io_73_DATA11    , hsma_io_74_DATA27   ,
			hsma_io_77_DATA12    , hsma_io_78_DATA28   ,
			hsma_io_79_DATA13    , hsma_io_80_DATA29   ,	
			hsma_io_83_DATA14    , hsma_io_84_DATA30   ,
			hsma_io_85_DATA15    , hsma_io_86_DATA31   ,
	
	output	hsma_out_d_101_BE_N[0]  		, hsma_out_d_102_TXE_N	,
			hsma_out_d_103_BE_N[1]  		, hsma_out_d_104_RXF_N	,
			hsma_out_d_107_BE_N[2]  		, hsma_out_d_108_SIWU_N	,
			hsma_out_d_109_BE_N[3]  		, hsma_out_d_110_WR_N	,
			hsma_out_d_113_GPIO_1_R_OOB   	, hsma_out_d_114_RD_N	,
			hsma_out_d_115_GPIO_0_W_OOB   	, hsma_out_d_116_OE_N	,
			hsma_out_d_119_RESET_N  		, 
			hsma_out_d_121_WAKEUP_N ; 
	
	
	
	