
package pkg_adc_defines ;


localparam 

ADC_WIDTH_DATA_IN 				= 12,
ADC_DESERIALIZATION_FACTOR 		= 8	,
ADC_WIDTH_DATA_DESER_OUT		= ADC_WIDTH_DATA_IN*ADC_DESERIALIZATION_FACTOR ,
ADC_WIDTH_DATA_FIFO_OUT			= 32,


	//FIFO_IN
			
	ADC_FIFO_IN_CNT_WORDS = 128,//Размером слова для FIFO является WIDTH_WRITE_DATA, т.е. он задается стороной записи 
	ADC_FIFO_IN_WIDTH_WRITE_DATA = ADC_WIDTH_DATA_DESER_OUT,
	ADC_FIFO_IN_WIDTH_READ_DATA = 32, //WIDTH_READ_DATA = 8и под него расчитывались размеры счетчиков
	ADC_FIFO_IN_COEFF_OTNOSHENIYA = ADC_FIFO_IN_WIDTH_WRITE_DATA/ADC_FIFO_IN_WIDTH_READ_DATA,
	ADC_FIFO_IN_WRITE_CNT =  $clog2(ADC_FIFO_IN_CNT_WORDS), // for this case = 10 
	ADC_FIFO_IN_READ_CNT = ( ADC_FIFO_IN_WIDTH_WRITE_DATA > ADC_FIFO_IN_WIDTH_READ_DATA ) ? ADC_FIFO_IN_WRITE_CNT + $clog2(ADC_FIFO_IN_COEFF_OTNOSHENIYA):  ADC_FIFO_IN_WRITE_CNT - $clog2(ADC_FIFO_IN_COEFF_OTNOSHENIYA),
	ADC_FIFO_IN_WIDTH_DELAY_PIPE = 4,

	VALUE_CNT_FIFO_IN_REDY_FOR_READ = ADC_FIFO_IN_CNT_WORDS/2,
	VALUE_CNT_FIFO_IN_END  = {(ADC_FIFO_IN_READ_CNT-1){1'b1}}


;



	
endpackage